`define module_name AHB_to_AHB_16_Bridge_Top
`define AHB_BUS_BASE_ADDR 32'hE8000000
`define AHB_SLAVE_ADDR_SIZE 4
`define AHB_SLAVE_1
